// create class with name usually corresponds to the specific task that you are performing. Acc to the architecture of our TB environment, each component will be built with the help of a class

class first;
  bit [2:0] data;  // declaring the data members of a class first
  bit [1:0] data2; // declaring the data members of a class first
endclass

// after finishing the declaration of a class, to utilize the class in the module, first create a handler
// by just creating a handler, you won't be able to access the class. The primary reason is that classes are dynamic objects, whereas the modules that we create are static objects. 
// STATIC VS DYNAMIC OBJECTS:  
//    when we perform a simulation from the start to the end of the simulation, "Module" object will be there. That is what we refer
//    to as static. Whereas when we consider a class, we may require it at some point during a simulation.
//    We do not keep that object alive for the entire simulation span. Instead, as and when required, we create an object, and once it serves its purpose, we delete it,
//    That is what we refer to as dynamic objects versus static objects, The modules defined here are static objects, 
//    so they are created at the start of a simulation and will stay till the end of the simulation, even if you do not utilize them during the entire simulation,


// Now let's try utilize a class inside a module, we can utilize in another class, package etc.,
module tb();
  first f;  // create a handler --> start with the class name, followed by a user-defined name for the handler. here f is the handler
            //  no memory is allocated to class and f points to a null
  first f2; // where we want to keep the original data as it is and utilize a copy of the original data for processing
 $display("Display1: Value of the data: %0d and data2 : %0d", f.data, f.data2); // if we use display without creating a constructor which means memory is not allocated, it gives NULL pointer error
  
  // all classes are dynamic. So we need to tell simulator when to allocate memory/ delete memory. So to allocate memory we create a object by adding a constructor
  //  we need to create a constructor that specifies when to create an object of a class. This is what we are doing to dynamically, when we need a class object, we create a constructor
  initial begin
    f = new();  // As soon as you add a constructor to the handler, memory is allocated for the class where the values of its data members will be stored, along with methods
                // Temporary data generated by the method will also be stored in that memory space,
                // Additionally, data members are initialized to their default values if the user does not initialize them. For a bit type, which represents a two-state value,
                // the default value is zero. For a four-state value (like reg), it will be initialized to x
    #1;
    $display("Display2:Value of the data: %0d and data2 : %0d", f.data, f.data2);

    // Now let's try to add values to the data memebers/properties
    // if we wan't to access Data members or methods of a class so, 'f' will act like a handler 
     f.data = 3'b101; 
     f.data2= 2'b10; 
     #1;
     $display("Display3: data: %0d and data2: %0d",f.data,f.data2);
    
     f = null ; // to deallocate the memory assigned to a class
     #1;
    $display("Display4: data: %0d and data2: %0d",f.data,f.data2);
  end
  
endmodule

// OUTPUT:
//KERNEL : fatal error : NULL POINTER ACCESS
//KERNEL : Display2: Value of the data: 0 and data2 0  // as data and data2 are bit datatype, default value is 0 // // if data and data2 are chnaged to reg datatype, default value is x
//kERNEL : Display3: Value of the data: 5 and data2 2  
//KERNEL : fatal error : NULL POINTER ACCESS

----------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
//////////////////////////////////// copying object by keeping original class ///////////////////////////////////
// where we want to keep the original data as it is and utilize a copy of the original data for processing
class first;
  int data;  // declaring the data members of a class first
  int data2; // declaring the data members of a class first
  function void display();
    $display("value of data: %0d, data2: %0d", data, data2);
  endfunction
endclass

module tb();
  first f1;  
  first f2; // where we want to keep the original data as it is and utilize a copy of the original data for processing
            // create another class veriable / handler
  first f3;
  initial begin
    f1 = new();  //// 1. call constructor for original class
    f1.data = 24; /// 2. Processing    
    f2 = new f1; //// 3. Create a copy from f1 to f2 . This creates a copy of the class. it copies all the data of f1 class into f2.
    $display("value of data member data from f1: %0d and data from f2: %0d",f1.data, f2.data); 
    f2.data = 32; //// Processing
    $display("value of data member data from f1: %0d and data from f2: %0d",f1.data, f2.data); 
    f3 = new();
    f1.data2 = 56;
    f3 = f1;   // create a copy  from f1 to f2
    f3.display();
    f1.display();
  end  
endmodule

// OUTPUT:
# KERNEL: value of data member data from f1: 24 and data from f2: 24
# KERNEL: value of data member data from f1: 24 and data from f2: 32
# KERNEL: value of data: 24, data2: 56
# KERNEL: value of data: 24, data2: 56

----------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
//////////////////////////////////// copying object - CUSTOM METHOD ///////////////////////////////////
//                  i. Add function inside class and Refer to add a constructor to the function name.   
//                   ii. So this will create an object, and once you have an object, you could just replace the data members of that object with the data of a claSS.  
//                  iii. In the testbench, you'll just call the custom method (function) that we have added, and this will return an object which we will store in the object where
class first;
  int data = 34;  // declaring the data members of a class first
  int data2; // declaring the data members of a class first
  function first copy();            // Add function inside class and Refer to add a constructor to the function name.
    copy = new();  /// 1. call constructor for original class to access datamembers
    copy.data = data;
    copy.data2 = data2;  
  endfunction
endclass

module tb();
  first f1, f2;  

  initial begin
    f1 = new();  //// 1. call constructor for original class
    f2 = new();
    f2 = f1.copy();        // In the testbench, you'll just call the custom method (function) that we have added, and this will return an object which we will store in the object 
     $display("value of data member data from f1: %0d and data from f2: %0d",f1.data, f2.data); 

  end  
endmodule

// OUTPUT:
//KERNEL : value of data member data from f1: 34 and data from f2: 34

----------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
//////////////////////////////////// copying object - SHALLOW COPY//////////////////////////////////////////////
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
----------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
//// here both original object and copied object has same handler
// get an independent copy of the data member but not an independent handler for both objects. that is refer to as a shallow copy. 
// that is why change in s2.f1.data will reflect the changes in s1.f1.data because both are pointing to same handler
// To have  both the original object and the copied object independent handlers, we use **"DEEP COPY"**

class first;
  int data =12;
endclass
class second;
    int data2 = 34;
    first f1;
    function new();
      f1 = new();
    endfunction
endclass

module tb;
  second s1, s2;
 initial begin 
   s1 = new();
   s1.data2= 45;
   s2 = new s1;
   $display("value of copied data2 : %0d",s2.data2); 
   s2.data2 = 78;
   $display("value of  data2in s1: %0d and s2: %0d", s1.data2, s2.data2);
   $display("value of  data in f1: %0d", s2.f1.data);
   s2.f1.data = 64;
   $display("value of  data in f1 from s1: %0d and from s2: %0d", s1.f1.data, s2.f1.data);
   
 end
endmodule

// OUTPUT:
# KERNEL: value of copied data2 : 45
# KERNEL: value of  data2in s1: 45 and s2: 78
# KERNEL: value of  data in f1: 12
# KERNEL: value of  data in f1: 64
# KERNEL: value of  data in f1 from s1: 64 and from s2: 64 // we get an independent copy of the data member but not an independent handler for both objects. that is refer to as a shallow copy
  
----------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
//////////////////////////////////// copying object - DEEP COPY//////////////////////////////////////////////
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
----------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
//// here both original object and copied object have different handler
// get an independent copy of the data member and independent copy of handler for both objects. that is refer to as a DEEP copy.
class first;
  int data =12;
  function first copy();           // Add function inside class and Refer to add a constructor to the function name.
    copy = new();  /// 1. call constructor for original class to access datamembers
    copy.data = data;
  endfunction
endclass
class second;
    int data2 = 34;
    first f1;
    function new();
      f1 = new();
    endfunction
  function second copy();             // Add function inside class and Refer to add a constructor to the function name.
    copy = new();  /// 1. call constructor for original class to access datamembers
    copy.data2 = data2;
    copy.f1 = f1.copy;
  endfunction
endclass

module tb;
  second s1, s2;
 initial begin 
   s1 = new();
   s2 = new();
   s1.data2= 45;
   s2 = s1.copy();
   $display("value of copied data2 : %0d",s2.data2); 
   s2.data2 = 78;
   $display("value of  data2in s1: %0d and s2: %0d", s1.data2, s2.data2);
   s2.f1.data = 64;
   $display("value of  data in f1 from s1: %0d and from s2: %0d", s1.f1.data, s2.f1.data);
   
 end
endmodule

// OUTPUT:
# KERNEL: value of copied data2 : 45
# KERNEL: value of  data2in s1: 45 and s2: 78
# KERNEL: value of  data in f1 from s1: 12 and from s2: 64
