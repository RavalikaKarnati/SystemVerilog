/////////////////////////////////////////////////////////////////////// TASK IN CLASS ///////////////////////////////////////////////////////////////////
