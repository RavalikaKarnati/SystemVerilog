// monitor
