
module tb;

class custom

endclass


endmodule
