module tb ();
  

endmodule
